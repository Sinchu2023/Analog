** sch_path: /foss/designs/Analog-Series/Day1/simulations/voltage_divider.sch
**.subckt voltage_divider
V1 n1 0 12v
R1 n1 vout 1k m=1
R2 vout 0 1k m=1
**** begin user architecture code

.dc v1 0 12 0.1

**** end user architecture code
**.ends
.end
